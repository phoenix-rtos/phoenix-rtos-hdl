-- UART 3
  constant CFG_UART3_ENABLE : integer := CONFIG_UART3_ENABLE;
  constant CFG_UART3_FIFO   : integer := CFG_UA3_FIFO;

