-- Xilinx MIG 7-Series
  constant CFG_MIG_7SERIES 	      : integer := CONFIG_MIG_ENABLE;
  constant CFG_MIG_7SERIES_MODEL  : integer := CONFIG_MIG_ENABLE;

