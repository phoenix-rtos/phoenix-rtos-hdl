-- LEON3 advanced interrupt controller
  constant CFG_IRQAMP_ENABLE: integer := CONFIG_IRQAMP_ENABLE;
-- LEON3 basic interrupt controller
  constant CFG_IRQ3_ENABLE  : integer := CONFIG_IRQ3_ENABLE;
  constant CFG_IRQ3_NSEC    : integer := CONFIG_IRQ3_NSEC;

